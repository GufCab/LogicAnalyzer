library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;
--library unisim;
--use unisim.vcomponents.all;

entity log_ctrl is
  generic (
    default_trig_chan : std_logic_vector(3 downto 0) := "0000";
  );
  port (
    
  );
end entity;
